module dac()